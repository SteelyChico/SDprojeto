`include "instruction_memory.sv"
`include "control_unit.sv"
`include "alu_control.sv"
`include "register_file.sv"
`include "alu.sv"
`include "data_memory.sv"
`include "sign_extend.sv"
`include "mips_processor.sv"
